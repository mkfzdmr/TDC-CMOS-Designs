* SPICE export by:  SEDIT 13.00
* Export time:      Thu Jan 31 22:56:52 2019
* Design:           Counter_TDC
* Cell:             schimit_trigger_2
* View:             view0
* Export as:        top-level cell
* Export mode:      hierarchical
* Exclude .model:   no
* Exclude .end:     no
* Expand paths:     yes
* Wrap lines:       no
* Root path:        C:\Users\makif\Google Drive\TEZ �ALI�MAM\�izim\Counter_TDC\Counter_TDC
* Exclude global pins:   no
* Control property name: SPICE

********* Simulation Settings - General section *********

********* Simulation Settings - Parameters and SPICE Options *********

*-------- Devices: SPICE.ORDER > 0 --------
MNMOS_1 N_1 In Gnd Out NMOS W=390n L=130n AS=351f PS=2.58u AD=351f PD=2.58u  
MNMOS_2 Out N_1 Gnd N_1 NMOS W=390n L=130n AS=351f PS=2.58u AD=351f PD=2.58u  
MPMOS_1 N_1 In Vdd Out PMOS W=390n L=130n AS=351f PS=2.58u AD=351f PD=2.58u  
MPMOS_2 Out N_1 Vdd N_1 PMOS W=390n L=130n AS=351f PS=2.58u AD=351f PD=2.58u  

********* Simulation Settings - Analysis section *********

********* Simulation Settings - Additional SPICE commands *********
VPower Vdd Gnd 1.4V
.include "C:\Users\makif\Google Drive\TEZ �ALI�MAM\�izim\�leri VLSI\VLSI_tech_files\130nm.md"
*.include "C:\Users\makif\Google Drive\TEZ �ALI�MAM\�izim\�leri VLSI\VLSI_tech_files\TSMC_0.18u_cmos.md"
*.include "C:\Users\makif\Google Drive\TEZ �ALI�MAM\�izim\�leri VLSI\VLSI_tech_files\SCN_0.25u_CMOS.md"
*.include "C:\Users\Hp\Google Drive\TEZ �ALI�MAM\�izim\�leri VLSI\VLSI_tech_files\130nm.md"
*.tran 0.01p 100p start=0


*VIn In Gnd BIT ({00001111} pw=5n lt=5n ht=5n on=3.3 off=0 rt=0.1n ft=0.1n delay=0)

VStart In 0 BIT ({0011111100} pw=10p lt=10p ht=10p on=1.4 off=0 rt=0.01p ft=0.01p delay=0)
*VStop Stop 0 BIT ({1110000000} pw=100n lt=100n ht=100n on=3.3 off=0 rt=0.01n ft=0.01n delay=0)

*VClock Clock 0 dc 0 PULSE (0 3.3V 0 0.001n 0.001n 0.6n 1.2n)
*VIn In 0 dc 0 PULSE (0 3.3 0 0.00000001n 0.00000001n 0.1n 0.02n)
*VIn In 0 dc 0 PULSE (0 3.3 0 0.1p 0.1p 10p 20p)

.tran 0.1p 100p start=0
.print tran   v(In,Gnd) v(Out,Gnd) 
*v(Start,Gnd) v(Stop,Gnd)
* v(INV_Q,Gnd)
.end

